package sequence_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "axi_lite_defines.svh"
    
    `include "axi_lite_seq_item.svh"
    `include "config_seq_item.svh"
    `include "axi_lite_sequence.svh"
    
endpackage: sequence_pkg