package analysis_components_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "axi_lite_defines.svh"

    import uvm_colors::*;
    import config_agent_pkg::*;
    import sequence_pkg::*;

    `include "config_checker.svh"
    `include "config_predictor.svh"
    `include "config_analysis_config.svh"
    
endpackage: analysis_components_pkg


