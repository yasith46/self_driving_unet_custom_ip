package config_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "axi_lite_defines.svh"

    import uvm_colors::*;
    import sequence_pkg::*;

    `include "config_agent_config.svh"
    `include "config_monitor.svh"
    `include "config_agent.svh"

endpackage: config_agent_pkg