package axi_lite_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "axi_lite_defines.svh"

    import uvm_colors::*;
    import sequence_pkg::*;

    `include "axi_lite_agent_config.svh"
    `include "axi_lite_monitor.svh"
    `include "axi_lite_slave_driver.svh"
    `include "axi_lite_agent.svh"

endpackage: axi_lite_agent_pkg