`define DATA_WIDTH 32