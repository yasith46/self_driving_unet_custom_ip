package axi_lite_test_pkg;

    import uvm_pkg::*;  
    `include "uvm_macros.svh"

    import axi_lite_agent_pkg::*;
    import env_pkg::*;
    import sequence_pkg::*;

    `include "axi_lite_defines.svh"
    `include    "axi_lite_test.svh"

endpackage: axi_lite_test_pkg